`include "const_def.v"

module ReOrderBuffer (

);

endmodule